library verilog;
use verilog.vl_types.all;
entity ascensor_vlg_vec_tst is
end ascensor_vlg_vec_tst;
