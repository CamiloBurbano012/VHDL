library verilog;
use verilog.vl_types.all;
entity puerta_vlg_vec_tst is
end puerta_vlg_vec_tst;
