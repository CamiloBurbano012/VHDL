library verilog;
use verilog.vl_types.all;
entity luces_vlg_check_tst is
    port(
        luz_cabina      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end luces_vlg_check_tst;
