library verilog;
use verilog.vl_types.all;
entity Panel_Fabrica_vlg_vec_tst is
end Panel_Fabrica_vlg_vec_tst;
