library verilog;
use verilog.vl_types.all;
entity Ascensor_vlg_vec_tst is
end Ascensor_vlg_vec_tst;
