library verilog;
use verilog.vl_types.all;
entity personas_vlg_vec_tst is
end personas_vlg_vec_tst;
