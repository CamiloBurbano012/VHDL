library verilog;
use verilog.vl_types.all;
entity Display_vlg_vec_tst is
end Display_vlg_vec_tst;
