library verilog;
use verilog.vl_types.all;
entity botones_vlg_vec_tst is
end botones_vlg_vec_tst;
