library verilog;
use verilog.vl_types.all;
entity motores_vlg_vec_tst is
end motores_vlg_vec_tst;
